`default_nettype none
`include "include/i2c.vh"
    
module i2c_tb;
endmodule

`default_nettype wire
